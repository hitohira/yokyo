module fdiv(
    input wire [31:0] x1,
    input wire [31:0] x2,
    output wire [31:0] y,
    input wire clk,
    input wire rstn);

    function [34:0] TDATA (
	input [9:0] MAL
    );
    begin
	casex(MAL)
        10'd0: TDATA = 35'b11111111110011111111100000000000100;
        10'd1: TDATA = 35'b11111111010011111110100000000100100;
        10'd2: TDATA = 35'b11111110110011111101100000001100100;
        10'd3: TDATA = 35'b11111110010011111100100000011000100;
        10'd4: TDATA = 35'b11111101110011111011100000101000100;
        10'd5: TDATA = 35'b11111101010011111010100000111100100;
        10'd6: TDATA = 35'b11111100110011111001100001010100100;
        10'd7: TDATA = 35'b11111100010011111000100001110000100;
        10'd8: TDATA = 35'b11111011110111110111101010001100010;
        10'd9: TDATA = 35'b11111011010111110110101010101111110;
        10'd10: TDATA = 35'b11111010110111110101101011010111010;
        10'd11: TDATA = 35'b11111010010111110100101100000010110;
        10'd12: TDATA = 35'b11111001110111110011101100110010010;
        10'd13: TDATA = 35'b11111001010111110010101101100101110;
        10'd14: TDATA = 35'b11111000111011110001110110010110001;
        10'd15: TDATA = 35'b11111000011011110000110111010001001;
        10'd16: TDATA = 35'b11110111111011101111111000010000001;
        10'd17: TDATA = 35'b11110111011011101110111001010011001;
        10'd18: TDATA = 35'b11110110111111101110000010010001000;
        10'd19: TDATA = 35'b11110110011111101101000011011011100;
        10'd20: TDATA = 35'b11110101111111101100000100101010000;
        10'd21: TDATA = 35'b11110101100011101011001101110010000;
        10'd22: TDATA = 35'b11110101000011101010001111001000000;
        10'd23: TDATA = 35'b11110100100011101001010000100010000;
        10'd24: TDATA = 35'b11110100000111101000011001110100000;
        10'd25: TDATA = 35'b11110011100111100111011011010101100;
        10'd26: TDATA = 35'b11110011000111100110011100111011000;
        10'd27: TDATA = 35'b11110010101011100101100110010111001;
        10'd28: TDATA = 35'b11110010001011100100101000000100001;
        10'd29: TDATA = 35'b11110001101111100011110001100110110;
        10'd30: TDATA = 35'b11110001001111100010110011011011010;
        10'd31: TDATA = 35'b11110000110011100001111101000100100;
        10'd32: TDATA = 35'b11110000010011100000111111000000100;
        10'd33: TDATA = 35'b11101111110011100000000001000000100;
        10'd34: TDATA = 35'b11101111010111011111001010110011110;
        10'd35: TDATA = 35'b11101110111011011110010100101010001;
        10'd36: TDATA = 35'b11101110011011011101010110110101001;
        10'd37: TDATA = 35'b11101101111111011100100000110010000;
        10'd38: TDATA = 35'b11101101011111011011100011000100100;
        10'd39: TDATA = 35'b11101101000011011010101101001000000;
        10'd40: TDATA = 35'b11101100100011011001101111100010000;
        10'd41: TDATA = 35'b11101100000111011000111001101100000;
        10'd42: TDATA = 35'b11101011101011011000000011111001001;
        10'd43: TDATA = 35'b11101011001011010111000110011110001;
        10'd44: TDATA = 35'b11101010101111010110010000110001110;
        10'd45: TDATA = 35'b11101010001111010101010011011110010;
        10'd46: TDATA = 35'b11101001110011010100011101111000100;
        10'd47: TDATA = 35'b11101001010111010011101000010101110;
        10'd48: TDATA = 35'b11101000111011010010110010110110001;
        10'd49: TDATA = 35'b11101000011011010001110101110001001;
        10'd50: TDATA = 35'b11100111111111010001000000011000000;
        10'd51: TDATA = 35'b11100111100011010000001011000010000;
        10'd52: TDATA = 35'b11100111000011001111001110001000000;
        10'd53: TDATA = 35'b11100110100111001110011000111000100;
        10'd54: TDATA = 35'b11100110001011001101100011101100001;
        10'd55: TDATA = 35'b11100101101111001100101110100010110;
        10'd56: TDATA = 35'b11100101010011001011111001011100100;
        10'd57: TDATA = 35'b11100100110011001010111100110100100;
        10'd58: TDATA = 35'b11100100010111001010000111110100110;
        10'd59: TDATA = 35'b11100011111011001001010010111000001;
        10'd60: TDATA = 35'b11100011011111001000011101111110100;
        10'd61: TDATA = 35'b11100011000011000111101001001000000;
        10'd62: TDATA = 35'b11100010100111000110110100010100100;
        10'd63: TDATA = 35'b11100010001011000101111111100100001;
        10'd64: TDATA = 35'b11100001101111000101001010110110110;
        10'd65: TDATA = 35'b11100001010011000100010110001100100;
        10'd66: TDATA = 35'b11100000110011000011011010000100100;
        10'd67: TDATA = 35'b11100000010111000010100101100000110;
        10'd68: TDATA = 35'b11011111111011000001110001000000001;
        10'd69: TDATA = 35'b11011111011111000000111100100010100;
        10'd70: TDATA = 35'b11011111000011000000001000001000000;
        10'd71: TDATA = 35'b11011110100110111111010011110000100;
        10'd72: TDATA = 35'b11011110001010111110011111011100001;
        10'd73: TDATA = 35'b11011101101110111101101011001010110;
        10'd74: TDATA = 35'b11011101010010111100110110111100100;
        10'd75: TDATA = 35'b11011100110110111100000010110001010;
        10'd76: TDATA = 35'b11011100011110111011010110000101100;
        10'd77: TDATA = 35'b11011100000010111010100010000000000;
        10'd78: TDATA = 35'b11011011100110111001101101111101100;
        10'd79: TDATA = 35'b11011011001010111000111001111110001;
        10'd80: TDATA = 35'b11011010101110111000000110000001110;
        10'd81: TDATA = 35'b11011010010010110111010010001000100;
        10'd82: TDATA = 35'b11011001110110110110011110010010010;
        10'd83: TDATA = 35'b11011001011010110101101010011111001;
        10'd84: TDATA = 35'b11011001000010110100111110001000000;
        10'd85: TDATA = 35'b11011000100110110100001010011010100;
        10'd86: TDATA = 35'b11011000001010110011010110110000001;
        10'd87: TDATA = 35'b11010111101110110010100011001000110;
        10'd88: TDATA = 35'b11010111010010110001101111100100100;
        10'd89: TDATA = 35'b11010110111010110001000011011010001;
        10'd90: TDATA = 35'b11010110011110110000001111111011100;
        10'd91: TDATA = 35'b11010110000010101111011100100000000;
        10'd92: TDATA = 35'b11010101100110101110101001000111100;
        10'd93: TDATA = 35'b11010101001110101101111101000111010;
        10'd94: TDATA = 35'b11010100110010101101001001110100100;
        10'd95: TDATA = 35'b11010100010110101100010110100100110;
        10'd96: TDATA = 35'b11010011111010101011100011011000001;
        10'd97: TDATA = 35'b11010011100010101010110111100010000;
        10'd98: TDATA = 35'b11010011000110101010000100011011000;
        10'd99: TDATA = 35'b11010010101010101001010001010111001;
        10'd100: TDATA = 35'b11010010010010101000100101101000100;
        10'd101: TDATA = 35'b11010001110110100111110010101010010;
        10'd102: TDATA = 35'b11010001011110100111000111000000100;
        10'd103: TDATA = 35'b11010001000010100110010100001000000;
        10'd104: TDATA = 35'b11010000100110100101100001010010100;
        10'd105: TDATA = 35'b11010000001110100100110101110000010;
        10'd106: TDATA = 35'b11001111110010100100000011000000100;
        10'd107: TDATA = 35'b11001111011010100011010111100011001;
        10'd108: TDATA = 35'b11001110111110100010100100111001000;
        10'd109: TDATA = 35'b11001110100110100001111001100000100;
        10'd110: TDATA = 35'b11001110001010100001000110111100001;
        10'd111: TDATA = 35'b11001101110010100000011011101000100;
        10'd112: TDATA = 35'b11001101010110011111101001001001110;
        10'd113: TDATA = 35'b11001100111110011110111101111011000;
        10'd114: TDATA = 35'b11001100100010011110001011100010000;
        10'd115: TDATA = 35'b11001100001010011101100000011000001;
        10'd116: TDATA = 35'b11001011101110011100101110000100110;
        10'd117: TDATA = 35'b11001011010110011100000010111111110;
        10'd118: TDATA = 35'b11001010111010011011010000110010001;
        10'd119: TDATA = 35'b11001010100010011010100101110010000;
        10'd120: TDATA = 35'b11001010000110011001110011101010000;
        10'd121: TDATA = 35'b11001001101110011001001000101110110;
        10'd122: TDATA = 35'b11001001010110011000011101110101110;
        10'd123: TDATA = 35'b11001000111010010111101011110110001;
        10'd124: TDATA = 35'b11001000100010010111000001000010000;
        10'd125: TDATA = 35'b11001000001010010110010110010000001;
        10'd126: TDATA = 35'b11000111101110010101100100011000110;
        10'd127: TDATA = 35'b11000111010110010100111001101011110;
        10'd128: TDATA = 35'b11000110111110010100001111000001000;
        10'd129: TDATA = 35'b11000110100010010011011101010010000;
        10'd130: TDATA = 35'b11000110001010010010110010101100001;
        10'd131: TDATA = 35'b11000101110010010010001000001000100;
        10'd132: TDATA = 35'b11000101010110010001010110100001110;
        10'd133: TDATA = 35'b11000100111110010000101100000011000;
        10'd134: TDATA = 35'b11000100100110010000000001100110100;
        10'd135: TDATA = 35'b11000100001110001111010111001100010;
        10'd136: TDATA = 35'b11000011110010001110100101110000100;
        10'd137: TDATA = 35'b11000011011010001101111011011011001;
        10'd138: TDATA = 35'b11000011000010001101010001001000000;
        10'd139: TDATA = 35'b11000010101010001100100110110111001;
        10'd140: TDATA = 35'b11000010010010001011111100101000100;
        10'd141: TDATA = 35'b11000001110110001011001011011010010;
        10'd142: TDATA = 35'b11000001011110001010100001010000100;
        10'd143: TDATA = 35'b11000001000110001001110111001001000;
        10'd144: TDATA = 35'b11000000101110001001001101000011110;
        10'd145: TDATA = 35'b11000000010110001000100011000000110;
        10'd146: TDATA = 35'b10111111111110000111111001000000000;
        10'd147: TDATA = 35'b10111111100110000111001111000001100;
        10'd148: TDATA = 35'b10111111001010000110011110000110001;
        10'd149: TDATA = 35'b10111110110010000101110100001100100;
        10'd150: TDATA = 35'b10111110011010000101001010010101001;
        10'd151: TDATA = 35'b10111110000010000100100000100000000;
        10'd152: TDATA = 35'b10111101101010000011110110101101001;
        10'd153: TDATA = 35'b10111101010010000011001100111100100;
        10'd154: TDATA = 35'b10111100111010000010100011001110001;
        10'd155: TDATA = 35'b10111100100010000001111001100010000;
        10'd156: TDATA = 35'b10111100001010000001001111111000001;
        10'd157: TDATA = 35'b10111011110010000000100110010000100;
        10'd158: TDATA = 35'b10111011011001111111111100101011001;
        10'd159: TDATA = 35'b10111011000001111111010011001000000;
        10'd160: TDATA = 35'b10111010101001111110101001100111001;
        10'd161: TDATA = 35'b10111010010001111110000000001000100;
        10'd162: TDATA = 35'b10111001111001111101010110101100001;
        10'd163: TDATA = 35'b10111001100001111100101101010010000;
        10'd164: TDATA = 35'b10111001001001111100000011111010001;
        10'd165: TDATA = 35'b10111000110001111011011010100100100;
        10'd166: TDATA = 35'b10111000011001111010110001010001001;
        10'd167: TDATA = 35'b10111000000001111010001000000000000;
        10'd168: TDATA = 35'b10110111101001111001011110110001001;
        10'd169: TDATA = 35'b10110111010101111000111100011011110;
        10'd170: TDATA = 35'b10110110111101111000010011010001000;
        10'd171: TDATA = 35'b10110110100101110111101010001000100;
        10'd172: TDATA = 35'b10110110001101110111000001000010010;
        10'd173: TDATA = 35'b10110101110101110110010111111110010;
        10'd174: TDATA = 35'b10110101011101110101101110111100100;
        10'd175: TDATA = 35'b10110101000101110101000101111101000;
        10'd176: TDATA = 35'b10110100110001110100100011110100100;
        10'd177: TDATA = 35'b10110100011001110011111010111001001;
        10'd178: TDATA = 35'b10110100000001110011010010000000000;
        10'd179: TDATA = 35'b10110011101001110010101001001001001;
        10'd180: TDATA = 35'b10110011010001110010000000010100100;
        10'd181: TDATA = 35'b10110010111101110001011110010101000;
        10'd182: TDATA = 35'b10110010100101110000110101100100100;
        10'd183: TDATA = 35'b10110010001101110000001100110110010;
        10'd184: TDATA = 35'b10110001110101101111100100001010010;
        10'd185: TDATA = 35'b10110001100001101111000010010010000;
        10'd186: TDATA = 35'b10110001001001101110011001101010001;
        10'd187: TDATA = 35'b10110000110001101101110001000100100;
        10'd188: TDATA = 35'b10110000011001101101001000100001001;
        10'd189: TDATA = 35'b10110000000101101100100110110000000;
        10'd190: TDATA = 35'b10101111101101101011111110010000110;
        10'd191: TDATA = 35'b10101111010101101011010101110011110;
        10'd192: TDATA = 35'b10101111000001101010110100001000000;
        10'd193: TDATA = 35'b10101110101001101010001011101111001;
        10'd194: TDATA = 35'b10101110010001101001100011011000100;
        10'd195: TDATA = 35'b10101101111101101001000001110010000;
        10'd196: TDATA = 35'b10101101100101101000011001011111100;
        10'd197: TDATA = 35'b10101101001101100111110001001111010;
        10'd198: TDATA = 35'b10101100111001100111001111101110001;
        10'd199: TDATA = 35'b10101100100001100110100111100010000;
        10'd200: TDATA = 35'b10101100001101100110000110000100010;
        10'd201: TDATA = 35'b10101011110101100101011101111100010;
        10'd202: TDATA = 35'b10101011011101100100110101110110100;
        10'd203: TDATA = 35'b10101011001001100100010100011110001;
        10'd204: TDATA = 35'b10101010110001100011101100011100100;
        10'd205: TDATA = 35'b10101010011101100011001011000111100;
        10'd206: TDATA = 35'b10101010000101100010100011001010000;
        10'd207: TDATA = 35'b10101001110001100010000001111000100;
        10'd208: TDATA = 35'b10101001011001100001011001111111001;
        10'd209: TDATA = 35'b10101001000101100000111000110001000;
        10'd210: TDATA = 35'b10101000101101100000010000111011110;
        10'd211: TDATA = 35'b10101000011001011111101111110001001;
        10'd212: TDATA = 35'b10101000000001011111001000000000000;
        10'd213: TDATA = 35'b10100111101101011110100110111000110;
        10'd214: TDATA = 35'b10100111010101011101111111001011110;
        10'd215: TDATA = 35'b10100111000001011101011110001000000;
        10'd216: TDATA = 35'b10100110101001011100110110011111001;
        10'd217: TDATA = 35'b10100110010101011100010101011110110;
        10'd218: TDATA = 35'b10100101111101011011101101111010000;
        10'd219: TDATA = 35'b10100101101001011011001100111101001;
        10'd220: TDATA = 35'b10100101010101011010101100000001110;
        10'd221: TDATA = 35'b10100100111101011010000100100011000;
        10'd222: TDATA = 35'b10100100101001011001100011101011001;
        10'd223: TDATA = 35'b10100100010001011000111100010000100;
        10'd224: TDATA = 35'b10100011111101011000011011011100000;
        10'd225: TDATA = 35'b10100011101001010111111010101001001;
        10'd226: TDATA = 35'b10100011010001010111010011010100100;
        10'd227: TDATA = 35'b10100010111101010110110010100101000;
        10'd228: TDATA = 35'b10100010100101010110001011010100100;
        10'd229: TDATA = 35'b10100010010001010101101010101000100;
        10'd230: TDATA = 35'b10100001111101010101001001111110000;
        10'd231: TDATA = 35'b10100001100101010100100010110011100;
        10'd232: TDATA = 35'b10100001010001010100000010001100100;
        10'd233: TDATA = 35'b10100000111101010011100001100111000;
        10'd234: TDATA = 35'b10100000101001010011000001000011001;
        10'd235: TDATA = 35'b10100000010001010010011010000000100;
        10'd236: TDATA = 35'b10011111111101010001111001100000000;
        10'd237: TDATA = 35'b10011111101001010001011001000001001;
        10'd238: TDATA = 35'b10011111010001010000110010000100100;
        10'd239: TDATA = 35'b10011110111101010000010001101001000;
        10'd240: TDATA = 35'b10011110101001001111110001001111001;
        10'd241: TDATA = 35'b10011110010101001111010000110110110;
        10'd242: TDATA = 35'b10011101111101001110101010000010000;
        10'd243: TDATA = 35'b10011101101001001110001001101101001;
        10'd244: TDATA = 35'b10011101010101001101101001011001110;
        10'd245: TDATA = 35'b10011101000001001101001001001000000;
        10'd246: TDATA = 35'b10011100101101001100101000110111110;
        10'd247: TDATA = 35'b10011100010101001100000010001100110;
        10'd248: TDATA = 35'b10011100000001001011100010000000000;
        10'd249: TDATA = 35'b10011011101101001011000001110100110;
        10'd250: TDATA = 35'b10011011011001001010100001101011001;
        10'd251: TDATA = 35'b10011011000101001010000001100011000;
        10'd252: TDATA = 35'b10011010110001001001100001011100100;
        10'd253: TDATA = 35'b10011010011001001000111010111101001;
        10'd254: TDATA = 35'b10011010000101001000011010111010000;
        10'd255: TDATA = 35'b10011001110001000111111010111000100;
        10'd256: TDATA = 35'b10011001011101000111011010111000100;
        10'd257: TDATA = 35'b10011001001001000110111010111010001;
        10'd258: TDATA = 35'b10011000110101000110011010111101010;
        10'd259: TDATA = 35'b10011000100001000101111011000010000;
        10'd260: TDATA = 35'b10011000001101000101011011001000010;
        10'd261: TDATA = 35'b10010111111001000100111011010000001;
        10'd262: TDATA = 35'b10010111100001000100010101000010000;
        10'd263: TDATA = 35'b10010111001101000011110101001101010;
        10'd264: TDATA = 35'b10010110111001000011010101011010001;
        10'd265: TDATA = 35'b10010110100101000010110101101000100;
        10'd266: TDATA = 35'b10010110010001000010010101111000100;
        10'd267: TDATA = 35'b10010101111101000001110110001010000;
        10'd268: TDATA = 35'b10010101101001000001010110011101001;
        10'd269: TDATA = 35'b10010101010101000000110110110001110;
        10'd270: TDATA = 35'b10010101000001000000010111001000000;
        10'd271: TDATA = 35'b10010100101100111111110111011111110;
        10'd272: TDATA = 35'b10010100011000111111010111111001001;
        10'd273: TDATA = 35'b10010100000100111110111000010100000;
        10'd274: TDATA = 35'b10010011110000111110011000110000100;
        10'd275: TDATA = 35'b10010011011100111101111001001110100;
        10'd276: TDATA = 35'b10010011001000111101011001101110001;
        10'd277: TDATA = 35'b10010010110100111100111010001111010;
        10'd278: TDATA = 35'b10010010100000111100011010110010000;
        10'd279: TDATA = 35'b10010010001100111011111011010110010;
        10'd280: TDATA = 35'b10010001111100111011100010001110000;
        10'd281: TDATA = 35'b10010001101000111011000010110101001;
        10'd282: TDATA = 35'b10010001010100111010100011011101110;
        10'd283: TDATA = 35'b10010001000000111010000100001000000;
        10'd284: TDATA = 35'b10010000101100111001100100110011110;
        10'd285: TDATA = 35'b10010000011000111001000101100001001;
        10'd286: TDATA = 35'b10010000000100111000100110010000000;
        10'd287: TDATA = 35'b10001111110000111000000111000000100;
        10'd288: TDATA = 35'b10001111011100110111100111110010100;
        10'd289: TDATA = 35'b10001111001000110111001000100110001;
        10'd290: TDATA = 35'b10001110111000110110101111101010001;
        10'd291: TDATA = 35'b10001110100100110110010000100000100;
        10'd292: TDATA = 35'b10001110010000110101110001011000100;
        10'd293: TDATA = 35'b10001101111100110101010010010010000;
        10'd294: TDATA = 35'b10001101101000110100110011001101001;
        10'd295: TDATA = 35'b10001101010100110100010100001001110;
        10'd296: TDATA = 35'b10001101000100110011111011010101000;
        10'd297: TDATA = 35'b10001100110000110011011100010100100;
        10'd298: TDATA = 35'b10001100011100110010111101010101100;
        10'd299: TDATA = 35'b10001100001000110010011110011000001;
        10'd300: TDATA = 35'b10001011110100110001111111011100010;
        10'd301: TDATA = 35'b10001011100100110001100110101101100;
        10'd302: TDATA = 35'b10001011010000110001000111110100100;
        10'd303: TDATA = 35'b10001010111100110000101000111101000;
        10'd304: TDATA = 35'b10001010101000110000001010000111001;
        10'd305: TDATA = 35'b10001010011000101111110001011101001;
        10'd306: TDATA = 35'b10001010000100101111010010101010000;
        10'd307: TDATA = 35'b10001001110000101110110011111000100;
        10'd308: TDATA = 35'b10001001011100101110010101001000100;
        10'd309: TDATA = 35'b10001001001100101101111100100011010;
        10'd310: TDATA = 35'b10001000111000101101011101110110001;
        10'd311: TDATA = 35'b10001000100100101100111111001010100;
        10'd312: TDATA = 35'b10001000010100101100100110101000110;
        10'd313: TDATA = 35'b10001000000000101100001000000000000;
        10'd314: TDATA = 35'b10000111101100101011101001011000110;
        10'd315: TDATA = 35'b10000111011000101011001010110011001;
        10'd316: TDATA = 35'b10000111001000101010110010010110001;
        10'd317: TDATA = 35'b10000110110100101010010011110011010;
        10'd318: TDATA = 35'b10000110100000101001110101010010000;
        10'd319: TDATA = 35'b10000110010000101001011100111000100;
        10'd320: TDATA = 35'b10000101111100101000111110011010000;
        10'd321: TDATA = 35'b10000101101100101000100110000010110;
        10'd322: TDATA = 35'b10000101011000101000000111100111001;
        10'd323: TDATA = 35'b10000101000100100111101001001101000;
        10'd324: TDATA = 35'b10000100110100100111010000111001010;
        10'd325: TDATA = 35'b10000100100000100110110010100010000;
        10'd326: TDATA = 35'b10000100001100100110010100001100010;
        10'd327: TDATA = 35'b10000011111100100101111011111100000;
        10'd328: TDATA = 35'b10000011101000100101011101101001001;
        10'd329: TDATA = 35'b10000011011000100101000101011011001;
        10'd330: TDATA = 35'b10000011000100100100100111001011000;
        10'd331: TDATA = 35'b10000010110100100100001110111111010;
        10'd332: TDATA = 35'b10000010100000100011110000110010000;
        10'd333: TDATA = 35'b10000010001100100011010010100110010;
        10'd334: TDATA = 35'b10000001111100100010111010011110000;
        10'd335: TDATA = 35'b10000001101000100010011100010101001;
        10'd336: TDATA = 35'b10000001011000100010000100001111001;
        10'd337: TDATA = 35'b10000001000100100001100110001001000;
        10'd338: TDATA = 35'b10000000110100100001001110000101010;
        10'd339: TDATA = 35'b10000000100000100000110000000010000;
        10'd340: TDATA = 35'b10000000010000100000011000000000100;
        10'd341: TDATA = 35'b01111111111100011111111010000000000;
        10'd342: TDATA = 35'b01111111101100011111100010000000110;
        10'd343: TDATA = 35'b01111111011000011111000100000011001;
        10'd344: TDATA = 35'b01111111001000011110101100000110001;
        10'd345: TDATA = 35'b01111110110100011110001110001011010;
        10'd346: TDATA = 35'b01111110100100011101110110010000100;
        10'd347: TDATA = 35'b01111110010000011101011000011000100;
        10'd348: TDATA = 35'b01111110000000011101000000100000000;
        10'd349: TDATA = 35'b01111101101100011100100010101010110;
        10'd350: TDATA = 35'b01111101011100011100001010110100100;
        10'd351: TDATA = 35'b01111101001100011011110010111111010;
        10'd352: TDATA = 35'b01111100111000011011010101001110001;
        10'd353: TDATA = 35'b01111100101000011010111101011011001;
        10'd354: TDATA = 35'b01111100010100011010011111101100110;
        10'd355: TDATA = 35'b01111100000100011010000111111100000;
        10'd356: TDATA = 35'b01111011110100011001110000001100010;
        10'd357: TDATA = 35'b01111011100000011001010010100010000;
        10'd358: TDATA = 35'b01111011010000011000111010110100100;
        10'd359: TDATA = 35'b01111010111100011000011101001101000;
        10'd360: TDATA = 35'b01111010101100011000000101100001110;
        10'd361: TDATA = 35'b01111010011100010111101101110111100;
        10'd362: TDATA = 35'b01111010001000010111010000010100001;
        10'd363: TDATA = 35'b01111001111000010110111000101100001;
        10'd364: TDATA = 35'b01111001100100010110011011001011100;
        10'd365: TDATA = 35'b01111001010100010110000011100101110;
        10'd366: TDATA = 35'b01111001000100010101101100000001000;
        10'd367: TDATA = 35'b01111000110000010101001110100100100;
        10'd368: TDATA = 35'b01111000100000010100110111000010000;
        10'd369: TDATA = 35'b01111000010000010100011111100000100;
        10'd370: TDATA = 35'b01110111111100010100000010001000000;
        10'd371: TDATA = 35'b01110111101100010011101010101000110;
        10'd372: TDATA = 35'b01110111011100010011010011001010100;
        10'd373: TDATA = 35'b01110111001100010010111011101101010;
        10'd374: TDATA = 35'b01110110111000010010011110011010001;
        10'd375: TDATA = 35'b01110110101000010010000110111111001;
        10'd376: TDATA = 35'b01110110011000010001101111100101001;
        10'd377: TDATA = 35'b01110110000100010001010010010110000;
        10'd378: TDATA = 35'b01110101110100010000111010111110010;
        10'd379: TDATA = 35'b01110101100100010000100011100111100;
        10'd380: TDATA = 35'b01110101010100010000001100010001110;
        10'd381: TDATA = 35'b01110101000000001111101111001000000;
        10'd382: TDATA = 35'b01110100110000001111010111110100100;
        10'd383: TDATA = 35'b01110100100000001111000000100010000;
        10'd384: TDATA = 35'b01110100010000001110101001010000100;
        10'd385: TDATA = 35'b01110011111100001110001100001100000;
        10'd386: TDATA = 35'b01110011101100001101110100111100110;
        10'd387: TDATA = 35'b01110011011100001101011101101110100;
        10'd388: TDATA = 35'b01110011001100001101000110100001010;
        10'd389: TDATA = 35'b01110010111100001100101111010101000;
        10'd390: TDATA = 35'b01110010101000001100010010010111001;
        10'd391: TDATA = 35'b01110010011000001011111011001101001;
        10'd392: TDATA = 35'b01110010001000001011100100000100001;
        10'd393: TDATA = 35'b01110001111000001011001100111100001;
        10'd394: TDATA = 35'b01110001101000001010110101110101001;
        10'd395: TDATA = 35'b01110001011000001010011110101111001;
        10'd396: TDATA = 35'b01110001000100001010000001111001000;
        10'd397: TDATA = 35'b01110000110100001001101010110101010;
        10'd398: TDATA = 35'b01110000100100001001010011110010100;
        10'd399: TDATA = 35'b01110000010100001000111100110000110;
        10'd400: TDATA = 35'b01110000000100001000100101110000000;
        10'd401: TDATA = 35'b01101111110100001000001110110000010;
        10'd402: TDATA = 35'b01101111100100000111110111110001100;
        10'd403: TDATA = 35'b01101111010000000111011011000100100;
        10'd404: TDATA = 35'b01101111000000000111000100001000000;
        10'd405: TDATA = 35'b01101110110000000110101101001100100;
        10'd406: TDATA = 35'b01101110100000000110010110010010000;
        10'd407: TDATA = 35'b01101110010000000101111111011000100;
        10'd408: TDATA = 35'b01101110000000000101101000100000000;
        10'd409: TDATA = 35'b01101101110000000101010001101000100;
        10'd410: TDATA = 35'b01101101100000000100111010110010000;
        10'd411: TDATA = 35'b01101101010000000100100011111100100;
        10'd412: TDATA = 35'b01101101000000000100001101001000000;
        10'd413: TDATA = 35'b01101100110000000011110110010100100;
        10'd414: TDATA = 35'b01101100011100000011011001110101100;
        10'd415: TDATA = 35'b01101100001100000011000011000100010;
        10'd416: TDATA = 35'b01101011111100000010101100010100000;
        10'd417: TDATA = 35'b01101011101100000010010101100100110;
        10'd418: TDATA = 35'b01101011011100000001111110110110100;
        10'd419: TDATA = 35'b01101011001100000001101000001001010;
        10'd420: TDATA = 35'b01101010111100000001010001011101000;
        10'd421: TDATA = 35'b01101010101100000000111010110001110;
        10'd422: TDATA = 35'b01101010011100000000100100000111100;
        10'd423: TDATA = 35'b01101010001100000000001101011110010;
        10'd424: TDATA = 35'b01101001111111111111101101101100000;
        10'd425: TDATA = 35'b01101001101111111111000000011101100;
        10'd426: TDATA = 35'b01101001011111111110010011010001000;
        10'd427: TDATA = 35'b01101001001111111101100110000110100;
        10'd428: TDATA = 35'b01101000111111111100111000111110000;
        10'd429: TDATA = 35'b01101000101111111100001011110111100;
        10'd430: TDATA = 35'b01101000011111111011011110110011000;
        10'd431: TDATA = 35'b01101000001111111010110001110000100;
        10'd432: TDATA = 35'b01100111111111111010000100110000000;
        10'd433: TDATA = 35'b01100111101111111001010111110001100;
        10'd434: TDATA = 35'b01100111100011111000110110000100000;
        10'd435: TDATA = 35'b01100111010011111000001001001001000;
        10'd436: TDATA = 35'b01100111000011110111011100010000000;
        10'd437: TDATA = 35'b01100110110011110110101111011001000;
        10'd438: TDATA = 35'b01100110100011110110000010100100000;
        10'd439: TDATA = 35'b01100110010011110101010101110001000;
        10'd440: TDATA = 35'b01100110000011110100101001000000000;
        10'd441: TDATA = 35'b01100101110011110011111100010001000;
        10'd442: TDATA = 35'b01100101100011110011001111100100000;
        10'd443: TDATA = 35'b01100101010011110010100010111001000;
        10'd444: TDATA = 35'b01100101000011110001110110010000000;
        10'd445: TDATA = 35'b01100100110011110001001001101001000;
        10'd446: TDATA = 35'b01100100100111110000101000001101000;
        10'd447: TDATA = 35'b01100100010111101111111011101001100;
        10'd448: TDATA = 35'b01100100000111101111001111001000000;
        10'd449: TDATA = 35'b01100011110111101110100010101000100;
        10'd450: TDATA = 35'b01100011100111101101110110001011000;
        10'd451: TDATA = 35'b01100011010111101101001001101111100;
        10'd452: TDATA = 35'b01100011000111101100011101010110000;
        10'd453: TDATA = 35'b01100010111011101011111100000100010;
        10'd454: TDATA = 35'b01100010101011101011001111101110010;
        10'd455: TDATA = 35'b01100010011011101010100011011010010;
        10'd456: TDATA = 35'b01100010001011101001110111001000010;
        10'd457: TDATA = 35'b01100001111011101001001010111000010;
        10'd458: TDATA = 35'b01100001101011101000011110101010010;
        10'd459: TDATA = 35'b01100001011111100111111101100001000;
        10'd460: TDATA = 35'b01100001001111100111010001010110100;
        10'd461: TDATA = 35'b01100000111111100110100101001110000;
        10'd462: TDATA = 35'b01100000101111100101111001000111100;
        10'd463: TDATA = 35'b01100000011111100101001101000011000;
        10'd464: TDATA = 35'b01100000010011100100101100000001000;
        10'd465: TDATA = 35'b01100000000011100100000000000000000;
        10'd466: TDATA = 35'b01011111110011100011010100000001000;
        10'd467: TDATA = 35'b01011111100011100010101000000100000;
        10'd468: TDATA = 35'b01011111010111100010000111000111100;
        10'd469: TDATA = 35'b01011111000111100001011011001110000;
        10'd470: TDATA = 35'b01011110110111100000101111010110100;
        10'd471: TDATA = 35'b01011110100111100000000011100001000;
        10'd472: TDATA = 35'b01011110010111011111010111101101100;
        10'd473: TDATA = 35'b01011110001011011110110110111000010;
        10'd474: TDATA = 35'b01011101111011011110001011001000010;
        10'd475: TDATA = 35'b01011101101011011101011111011010010;
        10'd476: TDATA = 35'b01011101011111011100111110101001000;
        10'd477: TDATA = 35'b01011101001111011100010010111110100;
        10'd478: TDATA = 35'b01011100111111011011100111010110000;
        10'd479: TDATA = 35'b01011100101111011010111011101111100;
        10'd480: TDATA = 35'b01011100100011011010011011000100000;
        10'd481: TDATA = 35'b01011100010011011001101111100001000;
        10'd482: TDATA = 35'b01011100000011011001000100000000000;
        10'd483: TDATA = 35'b01011011110111011000100011011000100;
        10'd484: TDATA = 35'b01011011100111010111110111111011000;
        10'd485: TDATA = 35'b01011011010111010111001100011111100;
        10'd486: TDATA = 35'b01011011001011010110101011111100010;
        10'd487: TDATA = 35'b01011010111011010110000000100100010;
        10'd488: TDATA = 35'b01011010101011010101010101001110010;
        10'd489: TDATA = 35'b01011010011111010100110100101111000;
        10'd490: TDATA = 35'b01011010001111010100001001011100100;
        10'd491: TDATA = 35'b01011001111111010011011110001100000;
        10'd492: TDATA = 35'b01011001110011010010111101110001000;
        10'd493: TDATA = 35'b01011001100011010010010010100100000;
        10'd494: TDATA = 35'b01011001010011010001100111011001000;
        10'd495: TDATA = 35'b01011001000111010001000111000010000;
        10'd496: TDATA = 35'b01011000110111010000011011111010100;
        10'd497: TDATA = 35'b01011000100111001111110000110101000;
        10'd498: TDATA = 35'b01011000011011001111010000100010010;
        10'd499: TDATA = 35'b01011000001011001110100101100000010;
        10'd500: TDATA = 35'b01010111111111001110000101010000000;
        10'd501: TDATA = 35'b01010111101111001101011010010001100;
        10'd502: TDATA = 35'b01010111011111001100101111010101000;
        10'd503: TDATA = 35'b01010111010011001100001111001001000;
        10'd504: TDATA = 35'b01010111000011001011100100010000000;
        10'd505: TDATA = 35'b01010110110111001011000100000110100;
        10'd506: TDATA = 35'b01010110100111001010011001010001000;
        10'd507: TDATA = 35'b01010110010111001001101110011101100;
        10'd508: TDATA = 35'b01010110001011001001001110011000010;
        10'd509: TDATA = 35'b01010101111011001000100011101000010;
        10'd510: TDATA = 35'b01010101101111001000000011100101100;
        10'd511: TDATA = 35'b01010101011111000111011000111001000;
        10'd512: TDATA = 35'b01010101010011000110111000111001000;
        10'd513: TDATA = 35'b01010101000011000110001110010000000;
        10'd514: TDATA = 35'b01010100110011000101100011101001000;
        10'd515: TDATA = 35'b01010100100111000101000011101101000;
        10'd516: TDATA = 35'b01010100010111000100011001001001100;
        10'd517: TDATA = 35'b01010100001011000011111001010000010;
        10'd518: TDATA = 35'b01010011111011000011001110110000010;
        10'd519: TDATA = 35'b01010011101111000010101110111001100;
        10'd520: TDATA = 35'b01010011011111000010000100011101000;
        10'd521: TDATA = 35'b01010011010011000001100100101001000;
        10'd522: TDATA = 35'b01010011000011000000111010010000000;
        10'd523: TDATA = 35'b01010010110111000000011010011110100;
        10'd524: TDATA = 35'b01010010100110111111110000001001000;
        10'd525: TDATA = 35'b01010010011010111111010000011010010;
        10'd526: TDATA = 35'b01010010001010111110100110001000010;
        10'd527: TDATA = 35'b01010001111110111110000110011100000;
        10'd528: TDATA = 35'b01010001101110111101011100001101100;
        10'd529: TDATA = 35'b01010001100010111100111100100100000;
        10'd530: TDATA = 35'b01010001010010111100010010011001000;
        10'd531: TDATA = 35'b01010001000110111011110010110010000;
        10'd532: TDATA = 35'b01010000110110111011001000101010100;
        10'd533: TDATA = 35'b01010000101010111010101001000110010;
        10'd534: TDATA = 35'b01010000011010111001111111000010010;
        10'd535: TDATA = 35'b01010000001110111001011111100000100;
        10'd536: TDATA = 35'b01010000000010111001000000000000000;
        10'd537: TDATA = 35'b01001111110010111000010110000001000;
        10'd538: TDATA = 35'b01001111100110110111110110100011000;
        10'd539: TDATA = 35'b01001111010110110111001100100111100;
        10'd540: TDATA = 35'b01001111001010110110101101001100010;
        10'd541: TDATA = 35'b01001110111010110110000011010100010;
        10'd542: TDATA = 35'b01001110101110110101100011111011100;
        10'd543: TDATA = 35'b01001110100010110101000100100100000;
        10'd544: TDATA = 35'b01001110010010110100011010110001000;
        10'd545: TDATA = 35'b01001110000110110011111011011100000;
        10'd546: TDATA = 35'b01001101110110110011010001101100100;
        10'd547: TDATA = 35'b01001101101010110010110010011010010;
        10'd548: TDATA = 35'b01001101011110110010010011001001000;
        10'd549: TDATA = 35'b01001101001110110001101001011110100;
        10'd550: TDATA = 35'b01001101000010110001001010010000000;
        10'd551: TDATA = 35'b01001100110010110000100000101001000;
        10'd552: TDATA = 35'b01001100100110110000000001011101000;
        10'd553: TDATA = 35'b01001100011010101111100010010010010;
        10'd554: TDATA = 35'b01001100001010101110111000110000010;
        10'd555: TDATA = 35'b01001011111110101110011001101000000;
        10'd556: TDATA = 35'b01001011110010101101111010100001000;
        10'd557: TDATA = 35'b01001011100010101101010001000100000;
        10'd558: TDATA = 35'b01001011010110101100110001111111100;
        10'd559: TDATA = 35'b01001011001010101100010010111100010;
        10'd560: TDATA = 35'b01001010111010101011101001100100010;
        10'd561: TDATA = 35'b01001010101110101011001010100011100;
        10'd562: TDATA = 35'b01001010011110101010100001001111000;
        10'd563: TDATA = 35'b01001010010010101010000010010001000;
        10'd564: TDATA = 35'b01001010000110101001100011010100000;
        10'd565: TDATA = 35'b01001001111010101001000100011000010;
        10'd566: TDATA = 35'b01001001101010101000011011001010010;
        10'd567: TDATA = 35'b01001001011110100111111100010001000;
        10'd568: TDATA = 35'b01001001010010100111011101011001000;
        10'd569: TDATA = 35'b01001001000010100110110100010000000;
        10'd570: TDATA = 35'b01001000110110100110010101011010100;
        10'd571: TDATA = 35'b01001000101010100101110110100110010;
        10'd572: TDATA = 35'b01001000011010100101001101100010010;
        10'd573: TDATA = 35'b01001000001110100100101110110000100;
        10'd574: TDATA = 35'b01001000000010100100010000000000000;
        10'd575: TDATA = 35'b01000111110110100011110001010000100;
        10'd576: TDATA = 35'b01000111100110100011001000010011000;
        10'd577: TDATA = 35'b01000111011010100010101001100110010;
        10'd578: TDATA = 35'b01000111001110100010001010111010100;
        10'd579: TDATA = 35'b01000110111110100001100010000010000;
        10'd580: TDATA = 35'b01000110110010100001000011011001000;
        10'd581: TDATA = 35'b01000110100110100000100100110001000;
        10'd582: TDATA = 35'b01000110011010100000000110001010010;
        10'd583: TDATA = 35'b01000110001010011111011101011000010;
        10'd584: TDATA = 35'b01000101111110011110111110110100000;
        10'd585: TDATA = 35'b01000101110010011110100000010001000;
        10'd586: TDATA = 35'b01000101100110011110000001101111000;
        10'd587: TDATA = 35'b01000101010110011101011001000011100;
        10'd588: TDATA = 35'b01000101001010011100111010100100010;
        10'd589: TDATA = 35'b01000100111110011100011100000110000;
        10'd590: TDATA = 35'b01000100110010011011111101101001000;
        10'd591: TDATA = 35'b01000100100110011011011111001101000;
        10'd592: TDATA = 35'b01000100010110011010110110101001100;
        10'd593: TDATA = 35'b01000100001010011010011000010000010;
        10'd594: TDATA = 35'b01000011111110011001111001111000000;
        10'd595: TDATA = 35'b01000011110010011001011011100001000;
        10'd596: TDATA = 35'b01000011100110011000111101001011000;
        10'd597: TDATA = 35'b01000011010110011000010100101111100;
        10'd598: TDATA = 35'b01000011001010010111110110011100010;
        10'd599: TDATA = 35'b01000010111110010111011000001010000;
        10'd600: TDATA = 35'b01000010110010010110111001111001000;
        10'd601: TDATA = 35'b01000010100110010110011011101001000;
        10'd602: TDATA = 35'b01000010010110010101110011010101100;
        10'd603: TDATA = 35'b01000010001010010101010101001000010;
        10'd604: TDATA = 35'b01000001111110010100110110111100000;
        10'd605: TDATA = 35'b01000001110010010100011000110001000;
        10'd606: TDATA = 35'b01000001100110010011111010100111000;
        10'd607: TDATA = 35'b01000001011010010011011100011110010;
        10'd608: TDATA = 35'b01000001001110010010111110010110100;
        10'd609: TDATA = 35'b01000000111110010010010110001110000;
        10'd610: TDATA = 35'b01000000110010010001111000001001000;
        10'd611: TDATA = 35'b01000000100110010001011010000101000;
        10'd612: TDATA = 35'b01000000011010010000111100000010010;
        10'd613: TDATA = 35'b01000000001110010000011110000000100;
        10'd614: TDATA = 35'b01000000000010010000000000000000000;
        10'd615: TDATA = 35'b00111111110110001111100010000000100;
        10'd616: TDATA = 35'b00111111100110001110111010000011000;
        10'd617: TDATA = 35'b00111111011010001110011100000110010;
        10'd618: TDATA = 35'b00111111001110001101111110001010100;
        10'd619: TDATA = 35'b00111111000010001101100000010000000;
        10'd620: TDATA = 35'b00111110110110001101000010010110100;
        10'd621: TDATA = 35'b00111110101010001100100100011110010;
        10'd622: TDATA = 35'b00111110011110001100000110100111000;
        10'd623: TDATA = 35'b00111110010010001011101000110001000;
        10'd624: TDATA = 35'b00111110000110001011001010111100000;
        10'd625: TDATA = 35'b00111101111010001010101101001000010;
        10'd626: TDATA = 35'b00111101101010001010000101011010010;
        10'd627: TDATA = 35'b00111101011110001001100111101001000;
        10'd628: TDATA = 35'b00111101010010001001001001111001000;
        10'd629: TDATA = 35'b00111101000110001000101100001010000;
        10'd630: TDATA = 35'b00111100111010001000001110011100010;
        10'd631: TDATA = 35'b00111100101110000111110000101111100;
        10'd632: TDATA = 35'b00111100100010000111010011000100000;
        10'd633: TDATA = 35'b00111100010110000110110101011001100;
        10'd634: TDATA = 35'b00111100001010000110010111110000010;
        10'd635: TDATA = 35'b00111011111110000101111010001000000;
        10'd636: TDATA = 35'b00111011110010000101011100100001000;
        10'd637: TDATA = 35'b00111011100110000100111110111011000;
        10'd638: TDATA = 35'b00111011011010000100100001010110010;
        10'd639: TDATA = 35'b00111011001110000100000011110010100;
        10'd640: TDATA = 35'b00111011000010000011100110010000000;
        10'd641: TDATA = 35'b00111010110110000011001000101110100;
        10'd642: TDATA = 35'b00111010101010000010101011001110010;
        10'd643: TDATA = 35'b00111010011110000010001101101111000;
        10'd644: TDATA = 35'b00111010010010000001110000010001000;
        10'd645: TDATA = 35'b00111010000110000001010010110100000;
        10'd646: TDATA = 35'b00111001111010000000110101011000010;
        10'd647: TDATA = 35'b00111001101110000000010111111101100;
        10'd648: TDATA = 35'b00111001100001111111111010100100000;
        10'd649: TDATA = 35'b00111001010101111111011101001011100;
        10'd650: TDATA = 35'b00111001001001111110111111110100010;
        10'd651: TDATA = 35'b00111000111101111110100010011110000;
        10'd652: TDATA = 35'b00111000110001111110000101001001000;
        10'd653: TDATA = 35'b00111000100101111101100111110101000;
        10'd654: TDATA = 35'b00111000011001111101001010100010010;
        10'd655: TDATA = 35'b00111000001101111100101101010000100;
        10'd656: TDATA = 35'b00111000000001111100010000000000000;
        10'd657: TDATA = 35'b00110111110101111011110010110000100;
        10'd658: TDATA = 35'b00110111101001111011010101100010010;
        10'd659: TDATA = 35'b00110111011101111010111000010101000;
        10'd660: TDATA = 35'b00110111010001111010011011001001000;
        10'd661: TDATA = 35'b00110111000101111001111101111110000;
        10'd662: TDATA = 35'b00110110111001111001100000110100010;
        10'd663: TDATA = 35'b00110110101101111001000011101011100;
        10'd664: TDATA = 35'b00110110100001111000100110100100000;
        10'd665: TDATA = 35'b00110110010101111000001001011101100;
        10'd666: TDATA = 35'b00110110001001110111101100011000010;
        10'd667: TDATA = 35'b00110101111101110111001111010100000;
        10'd668: TDATA = 35'b00110101110001110110110010010001000;
        10'd669: TDATA = 35'b00110101100101110110010101001111000;
        10'd670: TDATA = 35'b00110101011001110101111000001110010;
        10'd671: TDATA = 35'b00110101010001110101100100111001000;
        10'd672: TDATA = 35'b00110101000101110101000111111010000;
        10'd673: TDATA = 35'b00110100111001110100101010111100010;
        10'd674: TDATA = 35'b00110100101101110100001101111111100;
        10'd675: TDATA = 35'b00110100100001110011110001000100000;
        10'd676: TDATA = 35'b00110100010101110011010100001001100;
        10'd677: TDATA = 35'b00110100001001110010110111010000010;
        10'd678: TDATA = 35'b00110011111101110010011010011000000;
        10'd679: TDATA = 35'b00110011110001110001111101100001000;
        10'd680: TDATA = 35'b00110011100101110001100000101011000;
        10'd681: TDATA = 35'b00110011011101110001001101011101000;
        10'd682: TDATA = 35'b00110011010001110000110000101001000;
        10'd683: TDATA = 35'b00110011000101110000010011110110000;
        10'd684: TDATA = 35'b00110010111001101111110111000100010;
        10'd685: TDATA = 35'b00110010101101101111011010010011100;
        10'd686: TDATA = 35'b00110010100001101110111101100100000;
        10'd687: TDATA = 35'b00110010010101101110100000110101100;
        10'd688: TDATA = 35'b00110010001001101110000100001000010;
        10'd689: TDATA = 35'b00110010000001101101110001000000000;
        10'd690: TDATA = 35'b00110001110101101101010100010100100;
        10'd691: TDATA = 35'b00110001101001101100110111101010010;
        10'd692: TDATA = 35'b00110001011101101100011011000001000;
        10'd693: TDATA = 35'b00110001010001101011111110011001000;
        10'd694: TDATA = 35'b00110001000101101011100001110010000;
        10'd695: TDATA = 35'b00110000111101101011001110101110000;
        10'd696: TDATA = 35'b00110000110001101010110010001001000;
        10'd697: TDATA = 35'b00110000100101101010010101100101000;
        10'd698: TDATA = 35'b00110000011001101001111001000010010;
        10'd699: TDATA = 35'b00110000001101101001011100100000100;
        10'd700: TDATA = 35'b00110000000001101001000000000000000;
        10'd701: TDATA = 35'b00101111111001101000101101000000010;
        10'd702: TDATA = 35'b00101111101101101000010000100001100;
        10'd703: TDATA = 35'b00101111100001100111110100000100000;
        10'd704: TDATA = 35'b00101111010101100111010111100111100;
        10'd705: TDATA = 35'b00101111001001100110111011001100010;
        10'd706: TDATA = 35'b00101111000001100110101000010000000;
        10'd707: TDATA = 35'b00101110110101100110001011110110100;
        10'd708: TDATA = 35'b00101110101001100101101111011110010;
        10'd709: TDATA = 35'b00101110011101100101010011000111000;
        10'd710: TDATA = 35'b00101110010001100100110110110001000;
        10'd711: TDATA = 35'b00101110001001100100100011111000010;
        10'd712: TDATA = 35'b00101101111101100100000111100100000;
        10'd713: TDATA = 35'b00101101110001100011101011010001000;
        10'd714: TDATA = 35'b00101101100101100011001110111111000;
        10'd715: TDATA = 35'b00101101011001100010110010101110010;
        10'd716: TDATA = 35'b00101101010001100010011111111001000;
        10'd717: TDATA = 35'b00101101000101100010000011101010000;
        10'd718: TDATA = 35'b00101100111001100001100111011100010;
        10'd719: TDATA = 35'b00101100101101100001001011001111100;
        10'd720: TDATA = 35'b00101100100101100000111000011101000;
        10'd721: TDATA = 35'b00101100011001100000011100010010010;
        10'd722: TDATA = 35'b00101100001101100000000000001000100;
        10'd723: TDATA = 35'b00101100000001011111100100000000000;
        10'd724: TDATA = 35'b00101011111001011111010001010000010;
        10'd725: TDATA = 35'b00101011101101011110110101001001100;
        10'd726: TDATA = 35'b00101011100001011110011001000100000;
        10'd727: TDATA = 35'b00101011010101011101111100111111100;
        10'd728: TDATA = 35'b00101011001101011101101010010010100;
        10'd729: TDATA = 35'b00101011000001011101001110010000000;
        10'd730: TDATA = 35'b00101010110101011100110010001110100;
        10'd731: TDATA = 35'b00101010101001011100010110001110010;
        10'd732: TDATA = 35'b00101010100001011100000011100100000;
        10'd733: TDATA = 35'b00101010010101011011100111100101100;
        10'd734: TDATA = 35'b00101010001001011011001011101000010;
        10'd735: TDATA = 35'b00101010000001011010111001000000000;
        10'd736: TDATA = 35'b00101001110101011010011101000100100;
        10'd737: TDATA = 35'b00101001101001011010000001001010010;
        10'd738: TDATA = 35'b00101001011101011001100101010001000;
        10'd739: TDATA = 35'b00101001010101011001010010101011100;
        10'd740: TDATA = 35'b00101001001001011000110110110100010;
        10'd741: TDATA = 35'b00101000111101011000011010111110000;
        10'd742: TDATA = 35'b00101000110101011000001000011010100;
        10'd743: TDATA = 35'b00101000101001010111101100100110010;
        10'd744: TDATA = 35'b00101000011101010111010000110011000;
        10'd745: TDATA = 35'b00101000010101010110111110010001100;
        10'd746: TDATA = 35'b00101000001001010110100010100000010;
        10'd747: TDATA = 35'b00100111111101010110000110110000000;
        10'd748: TDATA = 35'b00100111110101010101110100010000100;
        10'd749: TDATA = 35'b00100111101001010101011000100010010;
        10'd750: TDATA = 35'b00100111011101010100111100110101000;
        10'd751: TDATA = 35'b00100111010101010100101010010111100;
        10'd752: TDATA = 35'b00100111001001010100001110101100010;
        10'd753: TDATA = 35'b00100110111101010011110011000010000;
        10'd754: TDATA = 35'b00100110110101010011100000100110100;
        10'd755: TDATA = 35'b00100110101001010011000100111110010;
        10'd756: TDATA = 35'b00100110011101010010101001010111000;
        10'd757: TDATA = 35'b00100110010101010010010110111101100;
        10'd758: TDATA = 35'b00100110001001010001111011011000010;
        10'd759: TDATA = 35'b00100101111101010001011111110100000;
        10'd760: TDATA = 35'b00100101110101010001001101011100100;
        10'd761: TDATA = 35'b00100101101001010000110001111010010;
        10'd762: TDATA = 35'b00100101100001010000011111100100000;
        10'd763: TDATA = 35'b00100101010101010000000100000011100;
        10'd764: TDATA = 35'b00100101001001001111101000100100010;
        10'd765: TDATA = 35'b00100101000001001111010110010000000;
        10'd766: TDATA = 35'b00100100110101001110111010110010100;
        10'd767: TDATA = 35'b00100100101001001110011111010110010;
        10'd768: TDATA = 35'b00100100100001001110001101000100000;
        10'd769: TDATA = 35'b00100100010101001101110001101001100;
        10'd770: TDATA = 35'b00100100001101001101011111011000100;
        10'd771: TDATA = 35'b00100100000001001101000100000000000;
        10'd772: TDATA = 35'b00100011110101001100101000101000100;
        10'd773: TDATA = 35'b00100011101101001100010110011001100;
        10'd774: TDATA = 35'b00100011100001001011111011000100000;
        10'd775: TDATA = 35'b00100011011001001011101000110110010;
        10'd776: TDATA = 35'b00100011001101001011001101100010100;
        10'd777: TDATA = 35'b00100011000001001010110010010000000;
        10'd778: TDATA = 35'b00100010111001001010100000000100010;
        10'd779: TDATA = 35'b00100010101101001010000100110011100;
        10'd780: TDATA = 35'b00100010100101001001110010101001000;
        10'd781: TDATA = 35'b00100010011001001001010111011010010;
        10'd782: TDATA = 35'b00100010010001001001000101010001000;
        10'd783: TDATA = 35'b00100010000101001000101010000100000;
        10'd784: TDATA = 35'b00100001111001001000001110111000010;
        10'd785: TDATA = 35'b00100001110001000111111100110001000;
        10'd786: TDATA = 35'b00100001100101000111100001100111000;
        10'd787: TDATA = 35'b00100001011101000111001111100001000;
        10'd788: TDATA = 35'b00100001010001000110110100011001000;
        10'd789: TDATA = 35'b00100001001001000110100010010100010;
        10'd790: TDATA = 35'b00100000111101000110000111001110000;
        10'd791: TDATA = 35'b00100000110101000101110101001010100;
        10'd792: TDATA = 35'b00100000101001000101011010000110010;
        10'd793: TDATA = 35'b00100000011101000100111111000011000;
        10'd794: TDATA = 35'b00100000010101000100101101000001100;
        10'd795: TDATA = 35'b00100000001001000100010010000000010;
        10'd796: TDATA = 35'b00100000000001000100000000000000000;
        10'd797: TDATA = 35'b00011111110101000011100101000000100;
        10'd798: TDATA = 35'b00011111101101000011010011000001100;
        10'd799: TDATA = 35'b00011111100001000010111000000100000;
        10'd800: TDATA = 35'b00011111011001000010100110000110010;
        10'd801: TDATA = 35'b00011111001101000010001011001010100;
        10'd802: TDATA = 35'b00011111000101000001111001001110000;
        10'd803: TDATA = 35'b00011110111001000001011110010100010;
        10'd804: TDATA = 35'b00011110110001000001001100011001000;
        10'd805: TDATA = 35'b00011110100101000000110001100001000;
        10'd806: TDATA = 35'b00011110011101000000011111100111000;
        10'd807: TDATA = 35'b00011110010001000000000100110001000;
        10'd808: TDATA = 35'b00011110001000111111110010111000010;
        10'd809: TDATA = 35'b00011101111100111111011000000100000;
        10'd810: TDATA = 35'b00011101110100111111000110001100100;
        10'd811: TDATA = 35'b00011101101000111110101011011010010;
        10'd812: TDATA = 35'b00011101100000111110011001100100000;
        10'd813: TDATA = 35'b00011101010100111101111110110011100;
        10'd814: TDATA = 35'b00011101001100111101101100111110100;
        10'd815: TDATA = 35'b00011101000000111101010010010000000;
        10'd816: TDATA = 35'b00011100111000111101000000011100010;
        10'd817: TDATA = 35'b00011100101100111100100101101111100;
        10'd818: TDATA = 35'b00011100100100111100010011111101000;
        10'd819: TDATA = 35'b00011100011000111011111001010010010;
        10'd820: TDATA = 35'b00011100010000111011100111100001000;
        10'd821: TDATA = 35'b00011100000100111011001100111000000;
        10'd822: TDATA = 35'b00011011111100111010111011001000000;
        10'd823: TDATA = 35'b00011011110100111010101001011000100;
        10'd824: TDATA = 35'b00011011101000111010001110110010010;
        10'd825: TDATA = 35'b00011011100000111001111101000100000;
        10'd826: TDATA = 35'b00011011010100111001100010011111100;
        10'd827: TDATA = 35'b00011011001100111001010000110010100;
        10'd828: TDATA = 35'b00011011000000111000110110010000000;
        10'd829: TDATA = 35'b00011010111000111000100100100100010;
        10'd830: TDATA = 35'b00011010101100111000001010000011100;
        10'd831: TDATA = 35'b00011010100100110111111000011001000;
        10'd832: TDATA = 35'b00011010011100110111100110101111000;
        10'd833: TDATA = 35'b00011010010000110111001100010001000;
        10'd834: TDATA = 35'b00011010001000110110111010101000010;
        10'd835: TDATA = 35'b00011001111100110110100000001100000;
        10'd836: TDATA = 35'b00011001110100110110001110100100100;
        10'd837: TDATA = 35'b00011001101000110101110100001010010;
        10'd838: TDATA = 35'b00011001100000110101100010100100000;
        10'd839: TDATA = 35'b00011001011000110101010000111110010;
        10'd840: TDATA = 35'b00011001001100110100110110100110100;
        10'd841: TDATA = 35'b00011001000100110100100101000010000;
        10'd842: TDATA = 35'b00011000111000110100001010101100010;
        10'd843: TDATA = 35'b00011000110000110011111001001001000;
        10'd844: TDATA = 35'b00011000100100110011011110110101000;
        10'd845: TDATA = 35'b00011000011100110011001101010011000;
        10'd846: TDATA = 35'b00011000010100110010111011110001100;
        10'd847: TDATA = 35'b00011000001000110010100001100000010;
        10'd848: TDATA = 35'b00011000000000110010010000000000000;
        10'd849: TDATA = 35'b00010111111000110001111110100000010;
        10'd850: TDATA = 35'b00010111101100110001100100010001100;
        10'd851: TDATA = 35'b00010111100100110001010010110011000;
        10'd852: TDATA = 35'b00010111011000110000111000100110010;
        10'd853: TDATA = 35'b00010111010000110000100111001001000;
        10'd854: TDATA = 35'b00010111001000110000010101101100010;
        10'd855: TDATA = 35'b00010110111100101111111011100010000;
        10'd856: TDATA = 35'b00010110110100101111101010000110100;
        10'd857: TDATA = 35'b00010110101000101111001111111110010;
        10'd858: TDATA = 35'b00010110100000101110111110100100000;
        10'd859: TDATA = 35'b00010110011000101110101101001010010;
        10'd860: TDATA = 35'b00010110001100101110010011000100100;
        10'd861: TDATA = 35'b00010110000100101110000001101100000;
        10'd862: TDATA = 35'b00010101111100101101110000010100000;
        10'd863: TDATA = 35'b00010101110000101101010110010001000;
        10'd864: TDATA = 35'b00010101101000101101000100111010010;
        10'd865: TDATA = 35'b00010101100000101100110011100100000;
        10'd866: TDATA = 35'b00010101010100101100011001100011100;
        10'd867: TDATA = 35'b00010101001100101100001000001110100;
        10'd868: TDATA = 35'b00010101000100101011110110111010000;
        10'd869: TDATA = 35'b00010100111000101011011100111100010;
        10'd870: TDATA = 35'b00010100110000101011001011101001000;
        10'd871: TDATA = 35'b00010100101000101010111010010110010;
        10'd872: TDATA = 35'b00010100011100101010100000011011000;
        10'd873: TDATA = 35'b00010100010100101010001111001001100;
        10'd874: TDATA = 35'b00010100001100101001111101111000100;
        10'd875: TDATA = 35'b00010100000000101001100100000000000;
        10'd876: TDATA = 35'b00010011111000101001010010110000010;
        10'd877: TDATA = 35'b00010011110000101001000001100001000;
        10'd878: TDATA = 35'b00010011100100101000100111101011000;
        10'd879: TDATA = 35'b00010011011100101000010110011101000;
        10'd880: TDATA = 35'b00010011010100101000000101001111100;
        10'd881: TDATA = 35'b00010011001000100111101011011100010;
        10'd882: TDATA = 35'b00010011000000100111011010010000000;
        10'd883: TDATA = 35'b00010010111000100111001001000100010;
        10'd884: TDATA = 35'b00010010101100100110101111010011100;
        10'd885: TDATA = 35'b00010010100100100110011110001001000;
        10'd886: TDATA = 35'b00010010011100100110001100111111000;
        10'd887: TDATA = 35'b00010010010000100101110011010001000;
        10'd888: TDATA = 35'b00010010001000100101100010001000010;
        10'd889: TDATA = 35'b00010010000000100101010001000000000;
        10'd890: TDATA = 35'b00010001111000100100111111111000010;
        10'd891: TDATA = 35'b00010001101100100100100110001101100;
        10'd892: TDATA = 35'b00010001100100100100010101000111000;
        10'd893: TDATA = 35'b00010001011100100100000100000001000;
        10'd894: TDATA = 35'b00010001010000100011101010011001000;
        10'd895: TDATA = 35'b00010001001000100011011001010100010;
        10'd896: TDATA = 35'b00010001000000100011001000010000000;
        10'd897: TDATA = 35'b00010000111000100010110111001100010;
        10'd898: TDATA = 35'b00010000101100100010011101100111100;
        10'd899: TDATA = 35'b00010000100100100010001100100101000;
        10'd900: TDATA = 35'b00010000011100100001111011100011000;
        10'd901: TDATA = 35'b00010000010100100001101010100001100;
        10'd902: TDATA = 35'b00010000001000100001010001000000010;
        10'd903: TDATA = 35'b00010000000000100001000000000000000;
        10'd904: TDATA = 35'b00001111111000100000101111000000010;
        10'd905: TDATA = 35'b00001111110000100000011110000001000;
        10'd906: TDATA = 35'b00001111100100100000000100100011000;
        10'd907: TDATA = 35'b00001111011100011111110011100101000;
        10'd908: TDATA = 35'b00001111010100011111100010100111100;
        10'd909: TDATA = 35'b00001111001100011111010001101010100;
        10'd910: TDATA = 35'b00001111000000011110111000010000000;
        10'd911: TDATA = 35'b00001110111000011110100111010100010;
        10'd912: TDATA = 35'b00001110110000011110010110011001000;
        10'd913: TDATA = 35'b00001110101000011110000101011110010;
        10'd914: TDATA = 35'b00001110011100011101101100000111000;
        10'd915: TDATA = 35'b00001110010100011101011011001101100;
        10'd916: TDATA = 35'b00001110001100011101001010010100100;
        10'd917: TDATA = 35'b00001110000100011100111001011100000;
        10'd918: TDATA = 35'b00001101111000011100100000001000010;
        10'd919: TDATA = 35'b00001101110000011100001111010001000;
        10'd920: TDATA = 35'b00001101101000011011111110011010010;
        10'd921: TDATA = 35'b00001101100000011011101101100100000;
        10'd922: TDATA = 35'b00001101011000011011011100101110010;
        10'd923: TDATA = 35'b00001101001100011011000011011110100;
        10'd924: TDATA = 35'b00001101000100011010110010101010000;
        10'd925: TDATA = 35'b00001100111100011010100001110110000;
        10'd926: TDATA = 35'b00001100110100011010010001000010100;
        10'd927: TDATA = 35'b00001100101100011010000000001111100;
        10'd928: TDATA = 35'b00001100100000011001100111000100000;
        10'd929: TDATA = 35'b00001100011000011001010110010010010;
        10'd930: TDATA = 35'b00001100010000011001000101100001000;
        10'd931: TDATA = 35'b00001100001000011000110100110000010;
        10'd932: TDATA = 35'b00001100000000011000100100000000000;
        10'd933: TDATA = 35'b00001011110100011000001010111000100;
        10'd934: TDATA = 35'b00001011101100010111111010001001100;
        10'd935: TDATA = 35'b00001011100100010111101001011011000;
        10'd936: TDATA = 35'b00001011011100010111011000101101000;
        10'd937: TDATA = 35'b00001011010100010111000111111111100;
        10'd938: TDATA = 35'b00001011001000010110101110111100010;
        10'd939: TDATA = 35'b00001011000000010110011110010000000;
        10'd940: TDATA = 35'b00001010111000010110001101100100010;
        10'd941: TDATA = 35'b00001010110000010101111100111001000;
        10'd942: TDATA = 35'b00001010101000010101101100001110010;
        10'd943: TDATA = 35'b00001010100000010101011011100100000;
        10'd944: TDATA = 35'b00001010010100010101000010100101100;
        10'd945: TDATA = 35'b00001010001100010100110001111100100;
        10'd946: TDATA = 35'b00001010000100010100100001010100000;
        10'd947: TDATA = 35'b00001001111100010100010000101100000;
        10'd948: TDATA = 35'b00001001110100010100000000000100100;
        10'd949: TDATA = 35'b00001001101100010011101111011101100;
        10'd950: TDATA = 35'b00001001100000010011010110100100000;
        10'd951: TDATA = 35'b00001001011000010011000101111110010;
        10'd952: TDATA = 35'b00001001010000010010110101011001000;
        10'd953: TDATA = 35'b00001001001000010010100100110100010;
        10'd954: TDATA = 35'b00001001000000010010010100010000000;
        10'd955: TDATA = 35'b00001000111000010010000011101100010;
        10'd956: TDATA = 35'b00001000110000010001110011001001000;
        10'd957: TDATA = 35'b00001000100100010001011010010101000;
        10'd958: TDATA = 35'b00001000011100010001001001110011000;
        10'd959: TDATA = 35'b00001000010100010000111001010001100;
        10'd960: TDATA = 35'b00001000001100010000101000110000100;
        10'd961: TDATA = 35'b00001000000100010000011000010000000;
        10'd962: TDATA = 35'b00000111111100010000000111110000000;
        10'd963: TDATA = 35'b00000111110100001111110111010000100;
        10'd964: TDATA = 35'b00000111101100001111100110110001100;
        10'd965: TDATA = 35'b00000111100000001111001110000100000;
        10'd966: TDATA = 35'b00000111011000001110111101100110010;
        10'd967: TDATA = 35'b00000111010000001110101101001001000;
        10'd968: TDATA = 35'b00000111001000001110011100101100010;
        10'd969: TDATA = 35'b00000111000000001110001100010000000;
        10'd970: TDATA = 35'b00000110111000001101111011110100010;
        10'd971: TDATA = 35'b00000110110000001101101011011001000;
        10'd972: TDATA = 35'b00000110101000001101011010111110010;
        10'd973: TDATA = 35'b00000110100000001101001010100100000;
        10'd974: TDATA = 35'b00000110010100001100110001111101100;
        10'd975: TDATA = 35'b00000110001100001100100001100100100;
        10'd976: TDATA = 35'b00000110000100001100010001001100000;
        10'd977: TDATA = 35'b00000101111100001100000000110100000;
        10'd978: TDATA = 35'b00000101110100001011110000011100100;
        10'd979: TDATA = 35'b00000101101100001011100000000101100;
        10'd980: TDATA = 35'b00000101100100001011001111101111000;
        10'd981: TDATA = 35'b00000101011100001010111111011001000;
        10'd982: TDATA = 35'b00000101010100001010101111000011100;
        10'd983: TDATA = 35'b00000101001100001010011110101110100;
        10'd984: TDATA = 35'b00000101000100001010001110011010000;
        10'd985: TDATA = 35'b00000100111000001001110101111100010;
        10'd986: TDATA = 35'b00000100110000001001100101101001000;
        10'd987: TDATA = 35'b00000100101000001001010101010110010;
        10'd988: TDATA = 35'b00000100100000001001000101000100000;
        10'd989: TDATA = 35'b00000100011000001000110100110010010;
        10'd990: TDATA = 35'b00000100010000001000100100100001000;
        10'd991: TDATA = 35'b00000100001000001000010100010000010;
        10'd992: TDATA = 35'b00000100000000001000000100000000000;
        10'd993: TDATA = 35'b00000011111000000111110011110000010;
        10'd994: TDATA = 35'b00000011110000000111100011100001000;
        10'd995: TDATA = 35'b00000011101000000111010011010010010;
        10'd996: TDATA = 35'b00000011100000000111000011000100000;
        10'd997: TDATA = 35'b00000011011000000110110010110110010;
        10'd998: TDATA = 35'b00000011010000000110100010101001000;
        10'd999: TDATA = 35'b00000011001000000110010010011100010;
        10'd1000: TDATA = 35'b00000011000000000110000010010000000;
        10'd1001: TDATA = 35'b00000010111000000101110010000100010;
        10'd1002: TDATA = 35'b00000010101100000101011001110011100;
        10'd1003: TDATA = 35'b00000010100100000101001001101001000;
        10'd1004: TDATA = 35'b00000010011100000100111001011111000;
        10'd1005: TDATA = 35'b00000010010100000100101001010101100;
        10'd1006: TDATA = 35'b00000010001100000100011001001100100;
        10'd1007: TDATA = 35'b00000010000100000100001001000100000;
        10'd1008: TDATA = 35'b00000001111100000011111000111100000;
        10'd1009: TDATA = 35'b00000001110100000011101000110100100;
        10'd1010: TDATA = 35'b00000001101100000011011000101101100;
        10'd1011: TDATA = 35'b00000001100100000011001000100111000;
        10'd1012: TDATA = 35'b00000001011100000010111000100001000;
        10'd1013: TDATA = 35'b00000001010100000010101000011011100;
        10'd1014: TDATA = 35'b00000001001100000010011000010110100;
        10'd1015: TDATA = 35'b00000001000100000010001000010010000;
        10'd1016: TDATA = 35'b00000000111100000001111000001110000;
        10'd1017: TDATA = 35'b00000000110100000001101000001010100;
        10'd1018: TDATA = 35'b00000000101100000001011000000111100;
        10'd1019: TDATA = 35'b00000000100100000001001000000101000;
        10'd1020: TDATA = 35'b00000000011100000000111000000011000;
        10'd1021: TDATA = 35'b00000000010100000000101000000001100;
        10'd1022: TDATA = 35'b00000000001100000000011000000000100;
        10'd1023: TDATA = 35'b00000000000100000000001000000000000;
        endcase
    end
    endfunction

    reg sy_reg1,sy_reg2;
    reg [7:0] ey0_reg1,ey1_reg1,ey0_reg2,ey1_reg2;
    reg [12:0] mx0_reg;
    reg [22:0] mx_reg1,mx_reg2,mix2_reg;
    reg [24:0] max02a_reg;

    // stage1
    wire sx,sy;
    wire [7:0] ex,ey;
    wire [22:0] mx,my;
    assign sx = x1[31];
    assign ex = x1[30:23];
    assign mx = x1[22:0];

    wire sa;
    wire [7:0] ea;
    wire [22:0] ma;
    assign sa = x2[31:31];
    assign ea = x2[30:23];
    assign ma = x2[22:0];

    assign sy = sx ^ sa;

    wire [9:0] mal;
    assign mal = x2[22:13];

    wire [34:0] tdata;
    assign tdata = TDATA(mal);
    
    wire [11:0] mx0;
    wire [22:0] mx02;
    assign mx0 = tdata[34:23];
    assign mx02 = tdata[22:0];

    wire [47:0] max02a;
    assign max02a = {1'b1,ma} * {1'b1,mx02};

    wire [8:0] eya0,eya1;
    assign eya0 = (ex == 0) ? 0: ex + 126;
    assign eya1 = (ex == 0) ? 0: ex + 127;

    wire [7:0] ey0,ey1;
    assign ey0 = (eya0 > ea) ? eya0 - ea: 0;
    assign ey1 = (eya1 > ea) ? eya1 - ea: 0;

    // stage2
    wire [22:0] max02;
    assign max02 = (max02a_reg[24]) ? max02a_reg[23:1]: max02a_reg[22:0];

    wire [24:0] mix2a;
    assign mix2a = {1'b1,mx0_reg,12'b0} - {2'b01,max02};

    wire [22:0] mix2;
    assign mix2 = mix2a[22:0];

    // stage3
    wire [47:0] mya;
    assign mya = {1'b1,mx_reg2} * {1'b1,mix2_reg};

    wire a;
    assign a = mya[47:47];
    assign my = (a) ? mya[46:24]: mya[45:23];
    assign ey = (a) ? ey1_reg2: ey0_reg2;

    assign y = {sy_reg2,ey,my};

    always @(posedge clk) begin
        // stage1
        sy_reg1 <= sy;
        mx_reg1 <= mx;
        mx0_reg <= mx0;
        max02a_reg <= max02a[47:23];
        ey0_reg1 <= ey0;
        ey1_reg1 <= ey1;

        // stage2
        sy_reg2 <= sy_reg1;
        mx_reg2 <= mx_reg1;
        mix2_reg <= mix2;
        ey0_reg2 <= ey0_reg1;
        ey1_reg2 <= ey1_reg1;

    end

    always @(negedge rstn) begin
       sy_reg1 <= 0;
       sy_reg2 <= 0; 
       ey0_reg1 <= 0;
       ey1_reg1 <= 0;
       ey0_reg2 <= 0;
       ey1_reg2 <= 0;
       mx0_reg <= 0;
       mx_reg1 <= 0;
       mx_reg2 <= 0;
       mix2_reg <= 0;
       max02a_reg <= 0;
    end

endmodule
